-- Copyright (C) 2021  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 21.1.0 Build 842 10/21/2021 SJ Lite Edition"
-- CREATED		"Sat Sep 14 15:19:44 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Block3 IS 
	PORT
	(
		T :  IN  STD_LOGIC;
		Clk :  IN  STD_LOGIC;
		Clear :  IN  STD_LOGIC;
		Q :  OUT  STD_LOGIC
	);
END Block3;

ARCHITECTURE bdf_type OF Block3 IS 



BEGIN 



PROCESS(Clk,Clear)
VARIABLE Q_synthesized_var : STD_LOGIC;
BEGIN
IF (Clear = '0') THEN
	Q_synthesized_var := '0';
ELSIF (RISING_EDGE(Clk)) THEN
	Q_synthesized_var := Q_synthesized_var XOR T;
END IF;
	Q <= Q_synthesized_var;
END PROCESS;


END bdf_type;